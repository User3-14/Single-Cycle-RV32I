-- Byte-offset controller - Store

library ieee;
use ieee.std_logic_1164.all;

entity Store_Control is
--	port (
--			
--		);
end entity;